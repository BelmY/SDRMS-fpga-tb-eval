
module cck (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
