
module rxpll (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
